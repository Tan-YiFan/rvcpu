module riscv_cpu_top (
  input         clock,
  input         reset,
  input         io_master_awready,
  output        io_master_awvalid,
  output [31:0] io_master_awaddr,
  output [2:0]  io_master_awprot,
  output        io_master_awid,
  output        io_master_awuser,
  output [7:0]  io_master_awlen,
  output [2:0]  io_master_awsize,
  output [1:0]  io_master_awburst,
  output        io_master_awlock,
  output [3:0]  io_master_awcache,
  output [3:0]  io_master_awqos,
  input         io_master_wready,
  output        io_master_wvalid,
  output [63:0] io_master_wdata,
  output [7:0]  io_master_wstrb,
  output        io_master_wlast,
  output        io_master_bready,
  input         io_master_bvalid,
  input  [1:0]  io_master_bresp,
  input         io_master_bid,
  input         io_master_buser,
  input         io_master_arready,
  output        io_master_arvalid,
  output [31:0] io_master_araddr,
  output [2:0]  io_master_arprot,
  output        io_master_arid,
  output        io_master_aruser,
  output [7:0]  io_master_arlen,
  output [2:0]  io_master_arsize,
  output [1:0]  io_master_arburst,
  output        io_master_arlock,
  output [3:0]  io_master_arcache,
  output [3:0]  io_master_arqos,
  output        io_master_rready,
  input         io_master_rvalid,
  input  [1:0]  io_master_rresp,
  input  [63:0] io_master_rdata,
  input         io_master_rlast,
  input         io_master_rid,
  input         io_master_ruser,
  input         io_interrupt
);
  /* riscv_cpu riscv_cpu (
    .clock(clock),
    .reset(reset),
    .io_mem_aw_ready(io_master_awready),
    .io_mem_aw_valid(io_master_awvalid),
    .io_mem_aw_bits_addr(io_master_awaddr),
    .io_mem_aw_bits_prot(io_master_awprot),
    .io_mem_aw_bits_id(io_master_awid),
    .io_mem_aw_bits_user(io_master_awuser),
    .io_mem_aw_bits_len(io_master_awlen),
    .io_mem_aw_bits_size(io_master_awsize),
    .io_mem_aw_bits_burst(io_master_awburst),
    .io_mem_aw_bits_lock(io_master_awlock),
    .io_mem_aw_bits_cache(io_master_awcache),
    .io_mem_aw_bits_qos(io_master_awqos),
    .io_mem_w_ready(io_master_wready),
    .io_mem_w_valid(io_master_wvalid),
    .io_mem_w_bits_data(io_master_wdata),
    .io_mem_w_bits_strb(io_master_wstrb),
    .io_mem_w_bits_last(io_master_wlast),
    .io_mem_b_ready(io_master_bready),
    .io_mem_b_valid(io_master_bvalid),
    .io_mem_b_bits_resp(io_master_bresp),
    .io_mem_b_bits_id(io_master_bid),
    .io_mem_b_bits_user(io_master_buser),
    .io_mem_ar_ready(io_master_arready),
    .io_mem_ar_valid(io_master_arvalid),
    .io_mem_ar_bits_addr(io_master_araddr),
    .io_mem_ar_bits_prot(io_master_arprot),
    .io_mem_ar_bits_id(io_master_arid),
    .io_mem_ar_bits_user(io_master_aruser),
    .io_mem_ar_bits_len(io_master_arlen),
    .io_mem_ar_bits_size(io_master_arsize),
    .io_mem_ar_bits_burst(io_master_arburst),
    .io_mem_ar_bits_lock(io_master_arlock),
    .io_mem_ar_bits_cache(io_master_arcache),
    .io_mem_ar_bits_qos(io_master_arqos),
    .io_mem_r_ready(io_master_rready),
    .io_mem_r_valid(io_master_rvalid),
    .io_mem_r_bits_resp(io_master_rresp),
    .io_mem_r_bits_data(io_master_rdata),
    .io_mem_r_bits_last(io_master_rlast),
    .io_mem_r_bits_id(io_master_rid),
    .io_mem_r_bits_user(io_master_ruser),
    .io_meip(io_interrupt)
  ); */

    mycpu_top mycpu_top (
    .clock(clock),
    .reset(reset),
    .awready(io_master_awready),
    .awvalid(io_master_awvalid),
    .awaddr(io_master_awaddr),
    .awprot(io_master_awprot),
    .awid(io_master_awid),
    .awuser(io_master_awuser),
    .awlen(io_master_awlen),
    .awsize(io_master_awsize),
    .awburst(io_master_awburst),
    .awlock(io_master_awlock),
    .awcache(io_master_awcache),
    .awqos(io_master_awqos),
    .wready(io_master_wready),
    .wvalid(io_master_wvalid),
    .wdata(io_master_wdata),
    .wstrb(io_master_wstrb),
    .wlast(io_master_wlast),
    .bready(io_master_bready),
    .bvalid(io_master_bvalid),
    .bresp(io_master_bresp),
    .bid(io_master_bid),
    .buser(io_master_buser),
    .arready(io_master_arready),
    .arvalid(io_master_arvalid),
    .araddr(io_master_araddr),
    .arprot(io_master_arprot),
    .arid(io_master_arid),
    .aruser(io_master_aruser),
    .arlen(io_master_arlen),
    .arsize(io_master_arsize),
    .arburst(io_master_arburst),
    .arlock(io_master_arlock),
    .arcache(io_master_arcache),
    .arqos(io_master_arqos),
    .rready(io_master_rready),
    .rvalid(io_master_rvalid),
    .rresp(io_master_rresp),
    .rdata(io_master_rdata),
    .rlast(io_master_rlast),
    .rid(io_master_rid),
    .ruser(io_master_ruser)
  );
endmodule
