`ifndef __EXCEPTION_PKG_SV
`define __EXCEPTION_PKG_SV



package exception_pkg;
	
endpackage

`endif
